module deco7segdec(

		input logic [3:0] D,
		output logic [6:0] SEG
	
);
//Este es el decodificador para las decenas
	always_comb begin
		case(D)
			4'b0000: SEG = 7'b1111111;
			4'b0001: SEG = 7'b1111001;
			4'b0010: SEG = 7'b0100100;
			4'b0011: SEG = 7'b0110000;
			4'b0100: SEG = 7'b0011001;
			4'b0101: SEG = 7'b0010010; 
			4'b0110: SEG = 7'b0000010;
			4'b0111: SEG = 7'b1111000;
			4'b1000: SEG = 7'b0000000;
			4'b1001: SEG = 7'b0011000;
			default: SEG = 7'b1111111;
		endcase
	end
endmodule
